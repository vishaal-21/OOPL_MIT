`timescale 1ns/1ns
`include "Q3.v"

module Q3_tb();
reg x1,x2,x3,x4,x5;
wire f;

Q3 P1(x1,x2,x3,x4,x5,f);
initial
begin
$dumpfile("Q3_tb.vcd");
$dumpvars(0, Q3_tb);
x1=0; x2=0; x3=0; x4=0; x5=0;
#20;
x1=0; x2=0; x3=0; x4=0; x5=1;
#20;
x1=0; x2=0; x3=0; x4=1; x5=0;
#20;
x1=0; x2=0; x3=0; x4=1; x5=1;
#20;
x1=0; x2=0; x3=1; x4=0; x5=0;
#20;
x1=0; x2=0; x3=1; x4=0; x5=1;
#20;
x1=0; x2=0; x3=1; x4=1; x5=0;
#20;
x1=0; x2=0; x3=1; x4=1; x5=1;
#20;
x1=0; x2=1; x3=0; x4=0; x5=0;
#20;
x1=0; x2=1; x3=0; x4=0; x5=1;
#20;
x1=0; x2=1; x3=0; x4=1; x5=0;
#20;
x1=0; x2=1; x3=0; x4=1; x5=1;
#20;
x1=0; x2=1; x3=1; x4=0; x5=0;
#20;
x1=0; x2=1; x3=1; x4=0; x5=1;
#20;
x1=0; x2=1; x3=1; x4=1; x5=0;
#20;
x1=0; x2=1; x3=1; x4=1; x5=1;
#20;
x1=1; x2=0; x3=0; x4=0; x5=0;
#20;
x1=1; x2=0; x3=0; x4=0; x5=1;
#20;
x1=1; x2=0; x3=0; x4=1; x5=0;
#20;
x1=1; x2=0; x3=0; x4=1; x5=1;
#20;
x1=1; x2=0; x3=1; x4=0; x5=0;
#20;
x1=1; x2=0; x3=1; x4=0; x5=1;
#20;
x1=1; x2=0; x3=1; x4=1; x5=0;
#20;
x1=1; x2=0; x3=1; x4=1; x5=1;
#20;
x1=1; x2=1; x3=0; x4=0; x5=0;
#20;
x1=1; x2=1; x3=0; x4=0; x5=1;
#20;
x1=1; x2=1; x3=0; x4=1; x5=0;
#20;
x1=1; x2=1; x3=0; x4=1; x5=1;
#20;
x1=1; x2=1; x3=1; x4=0; x5=0;
#20;
x1=1; x2=1; x3=1; x4=0; x5=1;
#20;
x1=1; x2=1; x3=1; x4=1; x5=0;
#20;
x1=1; x2=1; x3=1; x4=1; x5=1;
#20;
$display("Test complete");
end
endmodule
